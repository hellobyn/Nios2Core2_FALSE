// cpu2core.v

// Generated using ACDS version 14.1 186 at 2015.11.05.21:48:44

`timescale 1 ps / 1 ps
module cpu2core (
		input  wire        clk_clk,       //   clk.clk
		output wire        epcs_dclk,     //  epcs.dclk
		output wire        epcs_sce,      //      .sce
		output wire        epcs_sdo,      //      .sdo
		input  wire        epcs_data0,    //      .data0
		output wire [1:0]  pio0_export,   //  pio0.export
		input  wire        reset_reset_n, // reset.reset_n
		output wire [12:0] sdram_addr,    // sdram.addr
		output wire [1:0]  sdram_ba,      //      .ba
		output wire        sdram_cas_n,   //      .cas_n
		output wire        sdram_cke,     //      .cke
		output wire        sdram_cs_n,    //      .cs_n
		inout  wire [15:0] sdram_dq,      //      .dq
		output wire [1:0]  sdram_dqm,     //      .dqm
		output wire        sdram_ras_n,   //      .ras_n
		output wire        sdram_we_n     //      .we_n
	);

	wire  [31:0] cpu0_data_master_readdata;                                 // mm_interconnect_0:cpu0_data_master_readdata -> cpu0:d_readdata
	wire         cpu0_data_master_waitrequest;                              // mm_interconnect_0:cpu0_data_master_waitrequest -> cpu0:d_waitrequest
	wire         cpu0_data_master_debugaccess;                              // cpu0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu0_data_master_debugaccess
	wire  [26:0] cpu0_data_master_address;                                  // cpu0:d_address -> mm_interconnect_0:cpu0_data_master_address
	wire   [3:0] cpu0_data_master_byteenable;                               // cpu0:d_byteenable -> mm_interconnect_0:cpu0_data_master_byteenable
	wire         cpu0_data_master_read;                                     // cpu0:d_read -> mm_interconnect_0:cpu0_data_master_read
	wire         cpu0_data_master_write;                                    // cpu0:d_write -> mm_interconnect_0:cpu0_data_master_write
	wire  [31:0] cpu0_data_master_writedata;                                // cpu0:d_writedata -> mm_interconnect_0:cpu0_data_master_writedata
	wire  [31:0] cpu0_instruction_master_readdata;                          // mm_interconnect_0:cpu0_instruction_master_readdata -> cpu0:i_readdata
	wire         cpu0_instruction_master_waitrequest;                       // mm_interconnect_0:cpu0_instruction_master_waitrequest -> cpu0:i_waitrequest
	wire  [26:0] cpu0_instruction_master_address;                           // cpu0:i_address -> mm_interconnect_0:cpu0_instruction_master_address
	wire         cpu0_instruction_master_read;                              // cpu0:i_read -> mm_interconnect_0:cpu0_instruction_master_read
	wire         cpu0_instruction_master_readdatavalid;                     // mm_interconnect_0:cpu0_instruction_master_readdatavalid -> cpu0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_readdata;           // cpu0:debug_mem_slave_readdata -> mm_interconnect_0:cpu0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu0_debug_mem_slave_waitrequest;        // cpu0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu0_debug_mem_slave_debugaccess;        // mm_interconnect_0:cpu0_debug_mem_slave_debugaccess -> cpu0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu0_debug_mem_slave_address;            // mm_interconnect_0:cpu0_debug_mem_slave_address -> cpu0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu0_debug_mem_slave_read;               // mm_interconnect_0:cpu0_debug_mem_slave_read -> cpu0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu0_debug_mem_slave_byteenable;         // mm_interconnect_0:cpu0_debug_mem_slave_byteenable -> cpu0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu0_debug_mem_slave_write;              // mm_interconnect_0:cpu0_debug_mem_slave_write -> cpu0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu0_debug_mem_slave_writedata;          // mm_interconnect_0:cpu0_debug_mem_slave_writedata -> cpu0:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;       // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;         // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;          // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;             // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;            // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;        // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer0_s1_chipselect;                    // mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	wire  [15:0] mm_interconnect_0_timer0_s1_readdata;                      // timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer0_s1_address;                       // mm_interconnect_0:timer0_s1_address -> timer0:address
	wire         mm_interconnect_0_timer0_s1_write;                         // mm_interconnect_0:timer0_s1_write -> timer0:write_n
	wire  [15:0] mm_interconnect_0_timer0_s1_writedata;                     // mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	wire         mm_interconnect_0_pio0_s1_chipselect;                      // mm_interconnect_0:pio0_s1_chipselect -> pio0:chipselect
	wire  [31:0] mm_interconnect_0_pio0_s1_readdata;                        // pio0:readdata -> mm_interconnect_0:pio0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio0_s1_address;                         // mm_interconnect_0:pio0_s1_address -> pio0:address
	wire         mm_interconnect_0_pio0_s1_write;                           // mm_interconnect_0:pio0_s1_write -> pio0:write_n
	wire  [31:0] mm_interconnect_0_pio0_s1_writedata;                       // mm_interconnect_0:pio0_s1_writedata -> pio0:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // epcs:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu0_irq_irq;                                              // irq_mapper:sender_irq -> cpu0:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu0:reset_n, epcs:reset_n, irq_mapper:reset, mm_interconnect_0:cpu0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu0:reset_req, rst_translator:reset_req_in]
	wire         cpu0_debug_reset_request_reset;                            // cpu0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, pio0:reset_n, sdram:reset_n, sysid:reset_n, timer0:reset_n]

	cpu2core_cpu0 cpu0 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu0_data_master_read),                              //                          .read
		.d_readdata                          (cpu0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu0_data_master_write),                             //                          .write
		.d_writedata                         (cpu0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	cpu2core_epcs epcs (
		.clk           (clk_clk),                                             //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver1_irq),                            //               irq.irq
		.dclk          (epcs_dclk),                                           //          external.export
		.sce           (epcs_sce),                                            //                  .export
		.sdo           (epcs_sdo),                                            //                  .export
		.data0         (epcs_data0),                                          //                  .export
		.reset_req     (1'b0)                                                 //       (terminated)
	);

	cpu2core_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	cpu2core_pio0 pio0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_pio0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio0_s1_readdata),   //                    .readdata
		.out_port   (pio0_export)                           // external_connection.export
	);

	cpu2core_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	cpu2core_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	cpu2core_timer0 timer0 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                //   irq.irq
	);

	cpu2core_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                 (clk_clk),                                                   //                               clk_clk.clk
		.cpu0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                            //      cpu0_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu0_data_master_address                    (cpu0_data_master_address),                                  //                      cpu0_data_master.address
		.cpu0_data_master_waitrequest                (cpu0_data_master_waitrequest),                              //                                      .waitrequest
		.cpu0_data_master_byteenable                 (cpu0_data_master_byteenable),                               //                                      .byteenable
		.cpu0_data_master_read                       (cpu0_data_master_read),                                     //                                      .read
		.cpu0_data_master_readdata                   (cpu0_data_master_readdata),                                 //                                      .readdata
		.cpu0_data_master_write                      (cpu0_data_master_write),                                    //                                      .write
		.cpu0_data_master_writedata                  (cpu0_data_master_writedata),                                //                                      .writedata
		.cpu0_data_master_debugaccess                (cpu0_data_master_debugaccess),                              //                                      .debugaccess
		.cpu0_instruction_master_address             (cpu0_instruction_master_address),                           //               cpu0_instruction_master.address
		.cpu0_instruction_master_waitrequest         (cpu0_instruction_master_waitrequest),                       //                                      .waitrequest
		.cpu0_instruction_master_read                (cpu0_instruction_master_read),                              //                                      .read
		.cpu0_instruction_master_readdata            (cpu0_instruction_master_readdata),                          //                                      .readdata
		.cpu0_instruction_master_readdatavalid       (cpu0_instruction_master_readdatavalid),                     //                                      .readdatavalid
		.cpu0_debug_mem_slave_address                (mm_interconnect_0_cpu0_debug_mem_slave_address),            //                  cpu0_debug_mem_slave.address
		.cpu0_debug_mem_slave_write                  (mm_interconnect_0_cpu0_debug_mem_slave_write),              //                                      .write
		.cpu0_debug_mem_slave_read                   (mm_interconnect_0_cpu0_debug_mem_slave_read),               //                                      .read
		.cpu0_debug_mem_slave_readdata               (mm_interconnect_0_cpu0_debug_mem_slave_readdata),           //                                      .readdata
		.cpu0_debug_mem_slave_writedata              (mm_interconnect_0_cpu0_debug_mem_slave_writedata),          //                                      .writedata
		.cpu0_debug_mem_slave_byteenable             (mm_interconnect_0_cpu0_debug_mem_slave_byteenable),         //                                      .byteenable
		.cpu0_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu0_debug_mem_slave_waitrequest),        //                                      .waitrequest
		.cpu0_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu0_debug_mem_slave_debugaccess),        //                                      .debugaccess
		.epcs_epcs_control_port_address              (mm_interconnect_0_epcs_epcs_control_port_address),          //                epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                (mm_interconnect_0_epcs_epcs_control_port_write),            //                                      .write
		.epcs_epcs_control_port_read                 (mm_interconnect_0_epcs_epcs_control_port_read),             //                                      .read
		.epcs_epcs_control_port_readdata             (mm_interconnect_0_epcs_epcs_control_port_readdata),         //                                      .readdata
		.epcs_epcs_control_port_writedata            (mm_interconnect_0_epcs_epcs_control_port_writedata),        //                                      .writedata
		.epcs_epcs_control_port_chipselect           (mm_interconnect_0_epcs_epcs_control_port_chipselect),       //                                      .chipselect
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.pio0_s1_address                             (mm_interconnect_0_pio0_s1_address),                         //                               pio0_s1.address
		.pio0_s1_write                               (mm_interconnect_0_pio0_s1_write),                           //                                      .write
		.pio0_s1_readdata                            (mm_interconnect_0_pio0_s1_readdata),                        //                                      .readdata
		.pio0_s1_writedata                           (mm_interconnect_0_pio0_s1_writedata),                       //                                      .writedata
		.pio0_s1_chipselect                          (mm_interconnect_0_pio0_s1_chipselect),                      //                                      .chipselect
		.sdram_s1_address                            (mm_interconnect_0_sdram_s1_address),                        //                              sdram_s1.address
		.sdram_s1_write                              (mm_interconnect_0_sdram_s1_write),                          //                                      .write
		.sdram_s1_read                               (mm_interconnect_0_sdram_s1_read),                           //                                      .read
		.sdram_s1_readdata                           (mm_interconnect_0_sdram_s1_readdata),                       //                                      .readdata
		.sdram_s1_writedata                          (mm_interconnect_0_sdram_s1_writedata),                      //                                      .writedata
		.sdram_s1_byteenable                         (mm_interconnect_0_sdram_s1_byteenable),                     //                                      .byteenable
		.sdram_s1_readdatavalid                      (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                      .readdatavalid
		.sdram_s1_waitrequest                        (mm_interconnect_0_sdram_s1_waitrequest),                    //                                      .waitrequest
		.sdram_s1_chipselect                         (mm_interconnect_0_sdram_s1_chipselect),                     //                                      .chipselect
		.sysid_control_slave_address                 (mm_interconnect_0_sysid_control_slave_address),             //                   sysid_control_slave.address
		.sysid_control_slave_readdata                (mm_interconnect_0_sysid_control_slave_readdata),            //                                      .readdata
		.timer0_s1_address                           (mm_interconnect_0_timer0_s1_address),                       //                             timer0_s1.address
		.timer0_s1_write                             (mm_interconnect_0_timer0_s1_write),                         //                                      .write
		.timer0_s1_readdata                          (mm_interconnect_0_timer0_s1_readdata),                      //                                      .readdata
		.timer0_s1_writedata                         (mm_interconnect_0_timer0_s1_writedata),                     //                                      .writedata
		.timer0_s1_chipselect                        (mm_interconnect_0_timer0_s1_chipselect)                     //                                      .chipselect
	);

	cpu2core_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu0_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu0_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
