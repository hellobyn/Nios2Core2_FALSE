
module cpu2core (
	clk_clk,
	pio_0_export,
	pio_1_export,
	reset_reset_n);	

	input		clk_clk;
	output		pio_0_export;
	output		pio_1_export;
	input		reset_reset_n;
endmodule
