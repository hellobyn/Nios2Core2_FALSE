// cpu2core.v

// Generated using ACDS version 14.1 186 at 2015.11.03.21:03:28

`timescale 1 ps / 1 ps
module cpu2core (
		input  wire  clk_clk,       //   clk.clk
		output wire  pio_0_export,  // pio_0.export
		output wire  pio_1_export,  // pio_1.export
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_1_data_master_readdata;                                // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_waitrequest;                             // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire         cpu_1_data_master_debugaccess;                             // cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire  [16:0] cpu_1_data_master_address;                                 // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire   [3:0] cpu_1_data_master_byteenable;                              // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire         cpu_1_data_master_read;                                    // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire         cpu_1_data_master_write;                                   // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire  [31:0] cpu_1_data_master_writedata;                               // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire  [31:0] cpu_0_data_master_readdata;                                // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                             // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                             // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [16:0] cpu_0_data_master_address;                                 // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                              // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                    // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_write;                                   // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                               // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] cpu_0_instruction_master_readdata;                         // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                      // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [16:0] cpu_0_instruction_master_address;                          // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                             // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire  [31:0] cpu_1_instruction_master_readdata;                         // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire         cpu_1_instruction_master_waitrequest;                      // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire  [12:0] cpu_1_instruction_master_address;                          // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire         cpu_1_instruction_master_read;                             // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_readdata;          // cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest;       // cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess;       // mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1_debug_mem_slave_address;           // mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_read;              // mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1_debug_mem_slave_byteenable;        // mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_write;             // mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_writedata;         // mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_1_s1_chipselect;           // mm_interconnect_0:onchip_memory_1_s1_chipselect -> onchip_memory_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_1_s1_readdata;             // onchip_memory_1:readdata -> mm_interconnect_0:onchip_memory_1_s1_readdata
	wire   [7:0] mm_interconnect_0_onchip_memory_1_s1_address;              // mm_interconnect_0:onchip_memory_1_s1_address -> onchip_memory_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory_1_s1_byteenable;           // mm_interconnect_0:onchip_memory_1_s1_byteenable -> onchip_memory_1:byteenable
	wire         mm_interconnect_0_onchip_memory_1_s1_write;                // mm_interconnect_0:onchip_memory_1_s1_write -> onchip_memory_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory_1_s1_writedata;            // mm_interconnect_0:onchip_memory_1_s1_writedata -> onchip_memory_1:writedata
	wire         mm_interconnect_0_onchip_memory_1_s1_clken;                // mm_interconnect_0:onchip_memory_1_s1_clken -> onchip_memory_1:clken
	wire         mm_interconnect_0_pio_1_s1_chipselect;                     // mm_interconnect_0:pio_1_s1_chipselect -> pio_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;                       // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;                        // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_1_s1_write;                          // mm_interconnect_0:pio_1_s1_write -> pio_1:write_n
	wire  [31:0] mm_interconnect_0_pio_1_s1_writedata;                      // mm_interconnect_0:pio_1_s1_writedata -> pio_1:writedata
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;          // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;       // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;       // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;           // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_read;              // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;        // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_write;             // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;         // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_0_s1_chipselect;           // mm_interconnect_0:onchip_memory_0_s1_chipselect -> onchip_memory_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_0_s1_readdata;             // onchip_memory_0:readdata -> mm_interconnect_0:onchip_memory_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_0_s1_address;              // mm_interconnect_0:onchip_memory_0_s1_address -> onchip_memory_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory_0_s1_byteenable;           // mm_interconnect_0:onchip_memory_0_s1_byteenable -> onchip_memory_0:byteenable
	wire         mm_interconnect_0_onchip_memory_0_s1_write;                // mm_interconnect_0:onchip_memory_0_s1_write -> onchip_memory_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory_0_s1_writedata;            // mm_interconnect_0:onchip_memory_0_s1_writedata -> onchip_memory_0:writedata
	wire         mm_interconnect_0_onchip_memory_0_s1_clken;                // mm_interconnect_0:onchip_memory_0_s1_clken -> onchip_memory_0:clken
	wire         mm_interconnect_0_pio_0_s1_chipselect;                     // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                       // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                        // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                          // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                      // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver1_irq;                                  // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_0_irq_irq;                                             // irq_mapper:sender_irq -> cpu_0:irq
	wire  [31:0] cpu_1_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu_1:irq
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu_0:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, onchip_memory_0:reset, pio_0:reset_n, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu_0:reset_req, onchip_memory_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_0_debug_reset_request_reset;                           // cpu_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [cpu_1:reset_n, irq_mapper_001:reset, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, onchip_memory_1:reset, pio_1:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu_1:reset_req, onchip_memory_1:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_1_debug_reset_request_reset;                           // cpu_1:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, sysid:reset_n]

	cpu2core_cpu_0 cpu_0 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	cpu2core_cpu_1 cpu_1 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (cpu_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	cpu2core_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	cpu2core_onchip_memory_0 onchip_memory_0 (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)               //       .reset_req
	);

	cpu2core_onchip_memory_1 onchip_memory_1 (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)           //       .reset_req
	);

	cpu2core_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_export)                           // external_connection.export
	);

	cpu2core_pio_0 pio_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_1_s1_readdata),   //                    .readdata
		.out_port   (pio_1_export)                           // external_connection.export
	);

	cpu2core_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	cpu2core_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	cpu2core_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                 (clk_clk),                                                   //                               clk_clk.clk
		.cpu_0_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                            //     cpu_0_reset_reset_bridge_in_reset.reset
		.cpu_1_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                        //     cpu_1_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                   (cpu_0_data_master_address),                                 //                     cpu_0_data_master.address
		.cpu_0_data_master_waitrequest               (cpu_0_data_master_waitrequest),                             //                                      .waitrequest
		.cpu_0_data_master_byteenable                (cpu_0_data_master_byteenable),                              //                                      .byteenable
		.cpu_0_data_master_read                      (cpu_0_data_master_read),                                    //                                      .read
		.cpu_0_data_master_readdata                  (cpu_0_data_master_readdata),                                //                                      .readdata
		.cpu_0_data_master_write                     (cpu_0_data_master_write),                                   //                                      .write
		.cpu_0_data_master_writedata                 (cpu_0_data_master_writedata),                               //                                      .writedata
		.cpu_0_data_master_debugaccess               (cpu_0_data_master_debugaccess),                             //                                      .debugaccess
		.cpu_0_instruction_master_address            (cpu_0_instruction_master_address),                          //              cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest        (cpu_0_instruction_master_waitrequest),                      //                                      .waitrequest
		.cpu_0_instruction_master_read               (cpu_0_instruction_master_read),                             //                                      .read
		.cpu_0_instruction_master_readdata           (cpu_0_instruction_master_readdata),                         //                                      .readdata
		.cpu_1_data_master_address                   (cpu_1_data_master_address),                                 //                     cpu_1_data_master.address
		.cpu_1_data_master_waitrequest               (cpu_1_data_master_waitrequest),                             //                                      .waitrequest
		.cpu_1_data_master_byteenable                (cpu_1_data_master_byteenable),                              //                                      .byteenable
		.cpu_1_data_master_read                      (cpu_1_data_master_read),                                    //                                      .read
		.cpu_1_data_master_readdata                  (cpu_1_data_master_readdata),                                //                                      .readdata
		.cpu_1_data_master_write                     (cpu_1_data_master_write),                                   //                                      .write
		.cpu_1_data_master_writedata                 (cpu_1_data_master_writedata),                               //                                      .writedata
		.cpu_1_data_master_debugaccess               (cpu_1_data_master_debugaccess),                             //                                      .debugaccess
		.cpu_1_instruction_master_address            (cpu_1_instruction_master_address),                          //              cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest        (cpu_1_instruction_master_waitrequest),                      //                                      .waitrequest
		.cpu_1_instruction_master_read               (cpu_1_instruction_master_read),                             //                                      .read
		.cpu_1_instruction_master_readdata           (cpu_1_instruction_master_readdata),                         //                                      .readdata
		.cpu_0_debug_mem_slave_address               (mm_interconnect_0_cpu_0_debug_mem_slave_address),           //                 cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write                 (mm_interconnect_0_cpu_0_debug_mem_slave_write),             //                                      .write
		.cpu_0_debug_mem_slave_read                  (mm_interconnect_0_cpu_0_debug_mem_slave_read),              //                                      .read
		.cpu_0_debug_mem_slave_readdata              (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),          //                                      .readdata
		.cpu_0_debug_mem_slave_writedata             (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),         //                                      .writedata
		.cpu_0_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),        //                                      .byteenable
		.cpu_0_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),       //                                      .waitrequest
		.cpu_0_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),       //                                      .debugaccess
		.cpu_1_debug_mem_slave_address               (mm_interconnect_0_cpu_1_debug_mem_slave_address),           //                 cpu_1_debug_mem_slave.address
		.cpu_1_debug_mem_slave_write                 (mm_interconnect_0_cpu_1_debug_mem_slave_write),             //                                      .write
		.cpu_1_debug_mem_slave_read                  (mm_interconnect_0_cpu_1_debug_mem_slave_read),              //                                      .read
		.cpu_1_debug_mem_slave_readdata              (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),          //                                      .readdata
		.cpu_1_debug_mem_slave_writedata             (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),         //                                      .writedata
		.cpu_1_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),        //                                      .byteenable
		.cpu_1_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest),       //                                      .waitrequest
		.cpu_1_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess),       //                                      .debugaccess
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.onchip_memory_0_s1_address                  (mm_interconnect_0_onchip_memory_0_s1_address),              //                    onchip_memory_0_s1.address
		.onchip_memory_0_s1_write                    (mm_interconnect_0_onchip_memory_0_s1_write),                //                                      .write
		.onchip_memory_0_s1_readdata                 (mm_interconnect_0_onchip_memory_0_s1_readdata),             //                                      .readdata
		.onchip_memory_0_s1_writedata                (mm_interconnect_0_onchip_memory_0_s1_writedata),            //                                      .writedata
		.onchip_memory_0_s1_byteenable               (mm_interconnect_0_onchip_memory_0_s1_byteenable),           //                                      .byteenable
		.onchip_memory_0_s1_chipselect               (mm_interconnect_0_onchip_memory_0_s1_chipselect),           //                                      .chipselect
		.onchip_memory_0_s1_clken                    (mm_interconnect_0_onchip_memory_0_s1_clken),                //                                      .clken
		.onchip_memory_1_s1_address                  (mm_interconnect_0_onchip_memory_1_s1_address),              //                    onchip_memory_1_s1.address
		.onchip_memory_1_s1_write                    (mm_interconnect_0_onchip_memory_1_s1_write),                //                                      .write
		.onchip_memory_1_s1_readdata                 (mm_interconnect_0_onchip_memory_1_s1_readdata),             //                                      .readdata
		.onchip_memory_1_s1_writedata                (mm_interconnect_0_onchip_memory_1_s1_writedata),            //                                      .writedata
		.onchip_memory_1_s1_byteenable               (mm_interconnect_0_onchip_memory_1_s1_byteenable),           //                                      .byteenable
		.onchip_memory_1_s1_chipselect               (mm_interconnect_0_onchip_memory_1_s1_chipselect),           //                                      .chipselect
		.onchip_memory_1_s1_clken                    (mm_interconnect_0_onchip_memory_1_s1_clken),                //                                      .clken
		.pio_0_s1_address                            (mm_interconnect_0_pio_0_s1_address),                        //                              pio_0_s1.address
		.pio_0_s1_write                              (mm_interconnect_0_pio_0_s1_write),                          //                                      .write
		.pio_0_s1_readdata                           (mm_interconnect_0_pio_0_s1_readdata),                       //                                      .readdata
		.pio_0_s1_writedata                          (mm_interconnect_0_pio_0_s1_writedata),                      //                                      .writedata
		.pio_0_s1_chipselect                         (mm_interconnect_0_pio_0_s1_chipselect),                     //                                      .chipselect
		.pio_1_s1_address                            (mm_interconnect_0_pio_1_s1_address),                        //                              pio_1_s1.address
		.pio_1_s1_write                              (mm_interconnect_0_pio_1_s1_write),                          //                                      .write
		.pio_1_s1_readdata                           (mm_interconnect_0_pio_1_s1_readdata),                       //                                      .readdata
		.pio_1_s1_writedata                          (mm_interconnect_0_pio_1_s1_writedata),                      //                                      .writedata
		.pio_1_s1_chipselect                         (mm_interconnect_0_pio_1_s1_chipselect),                     //                                      .chipselect
		.sysid_control_slave_address                 (mm_interconnect_0_sysid_control_slave_address),             //                   sysid_control_slave.address
		.sysid_control_slave_readdata                (mm_interconnect_0_sysid_control_slave_readdata),            //                                      .readdata
		.timer_0_s1_address                          (mm_interconnect_0_timer_0_s1_address),                      //                            timer_0_s1.address
		.timer_0_s1_write                            (mm_interconnect_0_timer_0_s1_write),                        //                                      .write
		.timer_0_s1_readdata                         (mm_interconnect_0_timer_0_s1_readdata),                     //                                      .readdata
		.timer_0_s1_writedata                        (mm_interconnect_0_timer_0_s1_writedata),                    //                                      .writedata
		.timer_0_s1_chipselect                       (mm_interconnect_0_timer_0_s1_chipselect)                    //                                      .chipselect
	);

	cpu2core_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	cpu2core_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (cpu_1_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_0_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_1_debug_reset_request_reset),        // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
